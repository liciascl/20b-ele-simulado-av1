------------------------------
-- Elementos de Sistemas
-- Avaliacao Pratica 1
--
-- 10/2019
--
-- Questão 5
------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity q2 is
  port (
    x : in  STD_LOGIC_VECTOR(1 downto 0);
    y : in  STD_LOGIC_VECTOR(1 downto 0);
    z : out STD_LOGIC_VECTOR(3 downto 0));
end entity;

architecture  rtl OF q2 IS

begin


end architecture;
